------------------------------------------------
-- Switching element A_B
-- Acts as a router to link PEA and PEB
-- Lorenzo Lastrucci
------------------------------------------------
-- Entity Name       : AB_MUX
-- Architecture Name : STRUCT
------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use WORK.workpack.all;

entity AB_MUX is
 	port    (  X   :  in COMPLEX_ARRAY(0 to 31);
		   Y   : out COMPLEX_ARRAY(0 to 28);
		   SEL : in std_logic_vector(3 downto 0));
end AB_MUX;

architecture STRUCT of AB_MUX is
	constant O : COMPLEX := ((others=>'0'),(others=>'0'));
begin
	process(SEL,X)
	begin
		case SEL is
			when "0000" => 
				Y(0) <= X(0);
				Y(1) <= X(2);
				Y(2) <= X(4);
				Y(3) <= X(6);
				Y(4) <= X(8);
				Y(5) <= X(10);
				Y(6) <= X(12);
				Y(7) <= X(14);
				Y(8) <= X(16);
				Y(9) <= X(18);
				Y(10) <= X(20);
				Y(11) <= X(22);
				Y(12) <= X(24);
				Y(13) <= X(26);
				Y(14) <= X(28);
				Y(15) <= X(30);
				Y(16) <= O;
				Y(17) <= O;
				Y(18) <= O;
				Y(19) <= O;
				Y(20) <= O;
				Y(21) <= O;
				Y(22) <= O;
				Y(23) <= O;
				Y(24) <= O;
				Y(25) <= O;
				Y(26) <= O;
				Y(27) <= O;
				Y(28) <= O;
			when "0001" => 
				Y(0) <= X(1);
				Y(1) <= X(3);
				Y(2) <= X(5);
				Y(3) <= X(7);
				Y(4) <= X(9);
				Y(5) <= X(11);
				Y(6) <= X(13);
				Y(7) <= X(15);
				Y(8) <= X(17);
				Y(9) <= X(19);
				Y(10) <= X(21);
				Y(11) <= X(23);
				Y(12) <= X(25);
				Y(13) <= X(27);
				Y(14) <= X(29);
				Y(15) <= X(31);
				Y(16) <= O;
				Y(17) <= O;
				Y(18) <= O;
				Y(19) <= O;
				Y(20) <= O;
				Y(21) <= O;
				Y(22) <= O;
				Y(23) <= O;
				Y(24) <= O;
				Y(25) <= O;
				Y(26) <= O;
				Y(27) <= O;
				Y(28) <= O;
			when "1001" => 
				Y(0) <= O;
				Y(1) <= X(1);		--T32_1
				Y(2) <= X(3);		--T33_1
				Y(3) <= O;
				Y(4) <= X(9);		--T32_2
				Y(5) <= X(11);		--T33_2
				Y(6) <= O;
				Y(7) <= X(17);		--T32_3
				Y(8) <= X(19);		--T33_3
				Y(9) <= O;
				Y(10) <= X(25);		--T32_4
				Y(11) <= X(27);		--T33_4
				Y(12) <= O;
				Y(13) <= O;
				Y(14) <= O;
				Y(15) <= O;
				Y(16) <= X(6);		--T31_1
				Y(17) <= O;
				Y(18) <= X(14);		--T31_2
				Y(19) <= O;
				Y(20) <= O;
				Y(21) <= X(22);		--T31_3
				Y(22) <= O;
				Y(23) <= O;
				Y(24) <= X(30);		--T31_4
				Y(25) <= O;
				Y(26) <= O;
				Y(27) <= O;
				Y(28) <= O;
			when "1011" => 
				Y(0) <= O;
				Y(1) <= X(3);		--T55_1
				Y(2) <= O;
				Y(3) <= X(11);		--T56_1
				Y(4) <= O;
				Y(5) <= O;
				Y(6) <= O;
				Y(7) <= X(19);		--T55_2
				Y(8) <= O;
				Y(9) <= X(27);		--T56_2
				Y(10) <= O;
				Y(11) <= O;
				Y(12) <= O;
				Y(13) <= O;
				Y(14) <= O;
				Y(15) <= O;
				Y(16) <= X(6);		--T51_1
				Y(17) <= X(7);		--T58_1
				Y(18) <= X(22);		--T51_2
				Y(19) <= X(13);		--T59_1
				Y(20) <= O;
				Y(21) <= X(14);		--T53_1
				Y(22) <= X(29);		--T59_2
				Y(23) <= X(23);		--T58_2
				Y(24) <= X(30);		--T53_2
				Y(25) <= X(12);		--T52_1
				Y(26) <= X(1);		--T54_1
				Y(27) <= X(28);		--T52_2
				Y(28) <= X(17);		--T54_2
			when "1101" => 
				Y(0) <= X(1);		--T80_1
				Y(1) <= X(3);		--T84_1
				Y(2) <= X(5);		--T82_1
				Y(3) <= X(7);		--T86_1
				Y(4) <= X(9);		--T81_1
				Y(5) <= O;
				Y(6) <= O;
				Y(7) <= O;
				Y(8) <= X(17);		--T80_2
				Y(9) <= X(19);		--T84_2
				Y(10) <= X(21);		--T82_2
				Y(11) <= X(23);		--T86_2
				Y(12) <= X(25);		--T81_2
				Y(13) <= O;
				Y(14) <= O;
				Y(15) <= O;
				Y(16) <= O;
				Y(17) <= O;
				Y(18) <= O;
				Y(19) <= X(13);		--T83_1
				Y(20) <= X(11);		--T85_1
				Y(21) <= X(15);		--T87_1
				Y(22) <= X(29);		--T83_2
				Y(23) <= X(27);		--T85_2
				Y(24) <= X(31);		--T87_2
				Y(25) <= O;
				Y(26) <= O;
				Y(27) <= O;
				Y(28) <= O;
			when "1111" => 
				Y(0) <= X(1);		--T160
				Y(1) <= X(3);		--T168
				Y(2) <= X(5);		--T164
				Y(3) <= X(7);		--T1612
				Y(4) <= X(9);		--T161
				Y(5) <= O;
				Y(6) <= O;
				Y(7) <= O;
				Y(8) <= X(17);		--T162
				Y(9) <= O;
				Y(10) <= O;
				Y(11) <= O;
				Y(12) <= X(25);		--T163
				Y(13) <= O;
				Y(14) <= O;
				Y(15) <= O;
				Y(16) <= X(13);		--T165
				Y(17) <= X(21);		--T166
				Y(18) <= X(29);		--T167
				Y(19) <= X(11);		--T169
				Y(20) <= X(19);		--T1610
				Y(21) <= X(27);		--T1611
				Y(22) <= X(15);		--T1613
				Y(23) <= X(23);		--T1614
				Y(24) <= X(31);		--T1615
				Y(25) <= O;
				Y(26) <= O;
				Y(27) <= O;
				Y(28) <= O;
			when others => Y <= (others => O);
		end case;
	end process;
end STRUCT;








