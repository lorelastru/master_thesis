------------------------------------------------
-- Switching element B_C
-- Acts as a router to link PEB and PEC
-- Lorenzo Lastrucci
------------------------------------------------
-- Entity Name       : AB_MUX
-- Architecture Name : STRUCT
------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use WORK.workpack.all;

entity BC_MUX is
 	port    (  X   :  in COMPLEX_ARRAY(0 to 26);
		   Y   : out COMPLEX_ARRAY(0 to 19);
		   SEL : in std_logic_vector(3 downto 0));
end BC_MUX;

architecture STRUCT of BC_MUX is
	constant O : COMPLEX := ((others=>'0'),(others=>'0'));
begin
	process(SEL,X)
	begin
		case SEL is
			when "0000" => 		--radix_2
				Y(0) <= O;
				Y(1) <= O;
				Y(2) <= O;
				Y(3) <= O;
				Y(4) <= O;
				Y(5) <= O;
				Y(6) <= O;
				Y(7) <= O;
				Y(8) <= O;
				Y(9) <= O;
				Y(10) <= O;
				Y(11) <= O;
				Y(12) <= O;
				Y(13) <= O;
				Y(14) <= O;
				Y(15) <= O;
				Y(16) <= O;
				Y(17) <= O;
				Y(18) <= O;
				Y(19) <= O;
			when "0001" => 		--radix_4
				Y(0) <= O;
				Y(1) <= O;
				Y(2) <= O;
				Y(3) <= O;
				Y(4) <= O;
				Y(5) <= O;
				Y(6) <= O;
				Y(7) <= O;
				Y(8) <= O;
				Y(9) <= O;
				Y(10) <= O;
				Y(11) <= O;
				Y(12) <= O;
				Y(13) <= O;
				Y(14) <= O;
				Y(15) <= O;
				Y(16) <= O;
				Y(17) <= O;
				Y(18) <= O;
				Y(19) <= O;
			when "1001" => 		--radix_3
				Y(0) <= X(1);		--T32_1
				Y(1) <= X(4);		--T32_2
				Y(2) <= O;
				Y(3) <= O;
				Y(4) <= X(2);		--T33_1
				Y(5) <= X(16);		--M30_1	(T31_1)
				Y(6) <= O;
				Y(7) <= O;
				Y(8) <= X(5);		--T33_2
				Y(9) <= X(18);		--M30_2	(T31_2)
				Y(10) <= X(7);		--T32_3
				Y(11) <= X(10);		--T32_4
				Y(12) <= O;
				Y(13) <= O;
				Y(14) <= X(8);		--T33_3
				Y(15) <= X(21);		--M30_3	(T31_3)
				Y(16) <= O;
				Y(17) <= O;
				Y(18) <= X(11);		--T33_4
				Y(19) <= X(24);		--M30_4	(T31_4)
			when "1011" => 		--radix_5
				Y(0) <= X(25);		--T57_1
				Y(1) <= O;		
				Y(2) <= X(1);		--T55_1
				Y(3) <= X(17);		--M50_1	(T58_1)
				Y(4) <= X(17);		--M50_1	(T58_1)
				Y(5) <= X(3);		--T56_1
				Y(6) <= X(16);		--M53_1	(T51_1)
				Y(7) <= X(19);		--M52_1	(T59_1)
				Y(8) <= X(19);		--M52_1	(T59_1)
				Y(9) <= X(21);		--M51_1	(T53_1)
				Y(10) <= X(26);		--T57_2
				Y(11) <= O;		
				Y(12) <= X(7);		--T55_2
				Y(13) <= X(23);		--M50_2	(T58_2)
				Y(14) <= X(23);		--M50_2	(T58_2)
				Y(15) <= X(9);		--T56_2
				Y(16) <= X(18);		--M53_2 (T51_2)
				Y(17) <= X(22);		--M52_2	(T59_2)
				Y(18) <= X(22);		--M52_2	(T59_2)
				Y(19) <= X(24);		--M51_2	(T53_2)
			when "1101" => 		--radix_8
				Y(0) <= O;
				Y(1) <= O;
				Y(2) <= X(0);		--T80_1
				Y(3) <= X(4);		--T81_1
				Y(4) <= X(2);		--T82_1
				Y(5) <= X(19);		--M80_1 (T83_1)
				Y(6) <= X(1);		--T84_1
				Y(7) <= X(20);		--M81_1	(T85_1)
				Y(8) <= X(3);		--T86_1
				Y(9) <= X(21);		--M82_1	(T87_1)
				Y(10) <= O;
				Y(11) <= O;
				Y(12) <= X(8);		--T80_2	
				Y(13) <= X(12);		--T81_2
				Y(14) <= X(10);		--T82_2
				Y(15) <= X(22);		--M80_2	(T83_2)
				Y(16) <= X(9);		--T84_2
				Y(17) <= X(23);		--M81_2	(T85_2)
				Y(18) <= X(11);		--T86_2
				Y(19) <= X(24);		--M82_2	(T87_2)
			when "1111" => 		--radix_16
				Y(0) <= O;
				Y(1) <= O;
				Y(2) <= X(0);		--T160
				Y(3) <= X(8);		--T162
				Y(4) <= X(4);		--T161
				Y(5) <= X(12);		--T163
				Y(6) <= X(2);		--T164
				Y(7) <= X(17);		--M161	(T166)
				Y(8) <= X(16);		--M160	(T165)
				Y(9) <= X(18);		--M162	(T167)
				Y(10) <= O;
				Y(11) <= O;
				Y(12) <= X(1);		--T168
				Y(13) <= X(20);		--M164	(T1610)
				Y(14) <= X(19);		--M163	(T169)
				Y(15) <= X(21);		--M165	(T1611)
				Y(16) <= X(3);		--T1612
				Y(17) <= X(23);		--M167	(T1614)
				Y(18) <= X(22);		--M166	(T1613)
				Y(19) <= X(24);		--M168  (T1615)
			when others => Y <= (others => O);
		end case;
	end process;
end STRUCT;













